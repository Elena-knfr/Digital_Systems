module FA(a, b, cin, s, cout);
	input a, b, cin;
	output s, cout;
	
	assign s = cin ^ a ^ b;
	assign cout = (a & b) | (a & cin) | (b & cin);\
	
endmodule

	
